// =====================================
// MEM Stage (Memory Access)
// �t�d�G
//   - lw�GŪ��� memory[ALU_result]
//   - sw�G�g��� memory[ALU_result]
//   - ����T���ǻ��� MEM/WB
// =====================================

module MEM(
    input         clk,
    input         rst,

    // ===== EX/MEM pipeline inputs =====
    input         RegWrite_i,
    input         MemtoReg_i,
    input         MemRead_i,
    input         MemWrite_i,

    input  [31:0] ALU_result_i,   // memory address
    input  [31:0] rt_data_i,      // sw data
    input  [4:0]  dest_reg_i,     // �g�^���Ȧs���s��

    // ===== outputs to MEM/WB pipeline =====
    output        RegWrite_o,     // ���@����forwarding unit �i���o�䦳��ƭn�g�^, �@����MEM/WB
    output        MemtoReg_o,     // �~�򩹤U�Ǩ� WB ���q�� mux ���� �Ӧ۰O�����٬O ALU (ALU(0) / Memory(1, lw))
    output [31:0] read_data_o,    // lw data, �u�� MemRead=1 �ɤ~�|Ū
    output [31:0] ALU_result_o,   // bypass �� WB �H�� forwarding�ɻݭn
    output [4:0]  dest_reg_o      // to MEM/WB and forwarding unit
);

// =====================================
// DataMemory (lw / sw)
// =====================================
DataMemory DMEM(
    .clk        (clk),
    .MemRead_i  (MemRead_i),
    .MemWrite_i (MemWrite_i),
    .addr_i     (ALU_result_i),
    .write_data_i (rt_data_i),   // sw �����
    .read_data_o  (read_data_o)  // lw �����
);

// =====================================
// Pass signals to MEM/WB and forwarding unit
// =====================================
assign RegWrite_o   = RegWrite_i;       // to MEM/WB and forwarding unit
assign MemtoReg_o   = MemtoReg_i;       // to MEM/WB
assign ALU_result_o = ALU_result_i;     // to MEM/WB and forwarding unit and ALU mux
assign dest_reg_o   = dest_reg_i;       // to MEM/WB and forwarding unit

endmodule
