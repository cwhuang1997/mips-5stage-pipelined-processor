module EX_MEM(
    input clk, rst,

    // Control
    input RegWrite_i, MemtoReg_i, MemRead_i, MemWrite_i,
    // �O�_���\�⵲�G�g�^ Register File (R-type, lw, immmediate)
    // WB ���q�� mux ���� �Ӧ۰O�����٬O ALU (ALU(0) / Memory(1, lw))
    // �O����O�_�n���uŪ���v�ʧ@ (lw(1) / sw, R-type(0))
    // �O����O�_�n���u�g�J�v�ʧ@ (sw(1) / lw, R-type(0))

    // Data
    input [31:0] ALU_i,    // ALU result (�B�⵲�G, memory address)
    input [31:0] rt_i,     // ���F sw �n�g�J Data Memory ����� (�ĤG��mux�U������Output)
    input [4:0]  rd_i,     // �n�g�^���Ȧs���s��

    // Output
    output reg RegWrite_o, MemtoReg_o, MemRead_o, MemWrite_o,
    output reg [31:0] ALU_o,
    output reg [31:0] rt_o,
    output reg [4:0]  rd_o
);

always @(posedge clk or posedge rst) begin
    if (rst) begin
        {RegWrite_o, MemtoReg_o, MemRead_o, MemWrite_o} <= 0;
        ALU_o <= 0;
        rt_o  <= 0;
        rd_o  <= 0;
    end else begin
        RegWrite_o <= RegWrite_i;
        MemtoReg_o <= MemtoReg_i;
        MemRead_o  <= MemRead_i;
        MemWrite_o <= MemWrite_i;
    
        ALU_o <= ALU_i;
        rt_o  <= rt_i;
        rd_o  <= rd_i;
    end
end

endmodule
