// ===============================================
// Hazard Detection Unit
// �B�z lw-use hazard
// ===============================================
module Hazard_Detection_Unit(
    input        ID_EX_MemRead,    // EX ���q�����O�O�_�O lw
    input  [4:0] ID_EX_rt,         // lw ���ت��Ȧs�� (rt)

    input  [4:0] IF_ID_rs,         // �U�@�����O�� rs
    input  [4:0] IF_ID_rt,         // �U�@�����O�� rt

    output reg   PC_Write,         // PC_Write = 0 �� PC ���� ����s PC (�]�N�O�U�@�� clk��PC ����)
    output reg   IF_ID_Write,      // IF/ID Write = 0 �� IF/ID �Ȧs������s �O�����
    output reg   ID_EX_Flush,       // 1 �� ���J NOP�]�� EX �w 1 cycle�^


    input IF_ID_isBranch,
    input ID_EX_RegWrite,
    input [4:0] ID_EX_writeReg,
    input EX_MEM_RegWrite,
    input [4:0] EX_MEM_writeReg,
    input MEM_WB_RegWrite,
    input [4:0] MEM_WB_writeReg
);

always @(*) begin
    // �w�]���`�e�i�]�� stall�^
    PC_Write    = 1;
    IF_ID_Write = 1;
    ID_EX_Flush = 0;

    // ==========================
    // load-use hazard�G
    // lw $rt, XXX
    // �U�@�����O�p�G�ݭn rt �� forwarding �L�k�ѨM �� ���� stall
    // ==========================
    if (ID_EX_MemRead &&
       ((ID_EX_rt == IF_ID_rs) || (ID_EX_rt == IF_ID_rt))) begin    // �u�ˬd rt���S���ۦP(i.e., lw ���ت��Ȧs��) �t�@�ر��prs ��forwarding �ѨM

        PC_Write    = 0;   // PC ����]IF ���|���s���O�^
        IF_ID_Write = 0;   // IF/ID �Ȧs���O���]�קK�U�@���i�J EX�^
        ID_EX_Flush = 1;   // �b EX ���J bubble (NOP)
    end







    if (IF_ID_isBranch &&
        ID_EX_RegWrite &&
        (ID_EX_writeReg != 0) &&
        ((ID_EX_writeReg == IF_ID_rs) || (ID_EX_writeReg == IF_ID_rt)))
    begin
        PC_Write    = 0;
        IF_ID_Write = 0;
        ID_EX_Flush = 1;
    end

    if (IF_ID_isBranch &&
        EX_MEM_RegWrite &&
        (EX_MEM_writeReg != 0) &&
        ((EX_MEM_writeReg == IF_ID_rs) || (EX_MEM_writeReg == IF_ID_rt)))
    begin
        PC_Write    = 0;
        IF_ID_Write = 0;
        ID_EX_Flush = 1;
    end

    if (IF_ID_isBranch &&
        MEM_WB_RegWrite &&
        (MEM_WB_writeReg != 0) &&
        ((MEM_WB_writeReg == IF_ID_rs) || (MEM_WB_writeReg == IF_ID_rt)))
    begin
        PC_Write    = 0;
        IF_ID_Write = 0;
        ID_EX_Flush = 1;
    end




end

endmodule
