module IF_ID(
    input         clk,
    input         rst,              
    input         IF_ID_Write,      // hazard unit ����G1=��s, 0=�O�� (�Ω�load use hazard stalling)
    input  [31:0] instr_i,         // �q IF ���q�Ӫ����O
    input  [31:0] pc_i,            // �q IF ���q�Ӫ� PC+4
    output reg [31:0] instr_o,    // �� ID ���q�����O
    output reg [31:0] pc_o        // �� ID ���q�� PC+4
);

// �u���סGrst > IF_Flush > IF_ID_Write
always @(posedge clk or posedge rst) begin
    if (rst) begin
        instr_o <= 32'b0;
        pc_o    <= 32'b0;
    end 
    else if (IF_ID_Write) begin
        // Normal�G�S�� hazard �� pipeline ���`�y��
        instr_o <= instr_i;
        pc_o    <= pc_i;
    end
    // else: IF_ID_Write=0 �ɫO���{���ƭ�
end

endmodule
