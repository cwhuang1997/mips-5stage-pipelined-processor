// =====================================
// ID Stage (Instruction Decode)
// �t�d�G
//   1. Instruction Decode�]�� opcode ���ͱ���T���^
//   2. Register File �� Ū rs�Brt
//   3. Sign-Extend �� �ߧY���X�i�� 32-bit
//   4. Branch �P�_�]rs == rt�^
//   5. �N�Ҧ���ưe�� ID/EX pipeline register
// =====================================

module ID(
    input         clk,
    input         rst,

    // ===== �Ӧ� IF/ID Pipeline Register =====
    input  [31:0] instr_i,      // ���X�����O
    input  [31:0] pc_plus4_i,   // PC + 4�]�� branch �p��^

    // ===== �g�^���q�ݭn�g�^ RF =====
    input         WB_RegWrite_i, // (MEM/WB) RegWrite �H��
    // ���stage ���ʪ� RegWrite_in(1/0) ��F MEM/WB�� output �XWB_RegWrite_i(1/0)�Ǧ�Reg file
    input  [4:0]  WB_WriteAddr_i,// (MEM/WB) �g�^���ت��Ȧs�� (rd �� rt)
    input  [31:0] WB_WriteData_i,// (MEM/WB) �g�^�����

    // ===== ��X�� ID/EX Pipeline Register =====
    output        RegWrite_o,     // �O�_���\�g�^ Register File
    output        MemtoReg_o,     // WB mux�GALU(0) / Memory(1)
    output        MemRead_o,      // �O����Ū������ (lw=1 / ��L=0)
    output        MemWrite_o,     // �O����g�J���� (sw=1 / ��L=0)
    output [1:0]  ALUOp_o,        // ALU �B��X
    output        ALUSrc_o,       // ALU �ĤG�B�⤸�G�H�s��(0) / �ߧY��(1)

    output [31:0] rs_data_o,      // rs �H�s�����
    output [31:0] rt_data_o,      // rt �H�s�����
    output [31:0] imm_o,          // �Ÿ��X�i�᪺�ߧY��
    output [5:0]  funct_o,        // funct field�]�Ω� ALU Control�^

    output [4:0]  rs_addr_o,      // rs ��}
    output [4:0]  rt_addr_o,      // rt ��}
    output [4:0]  rd_addr_o,      // rd ��}

    // ===== BEQ  =====
    output        Branch_o, 
    output        Zero_o,              // rs == rt ?
    output [31:0] branch_target_o      // PC + 4 + (imm << 2)
);

wire [5:0] opcode  = instr_i[31:26];
wire [4:0] rs      = instr_i[25:21];
wire [4:0] rt      = instr_i[20:16];
wire [4:0] rd      = instr_i[15:11];
wire [5:0] funct   = instr_i[5:0];
wire [15:0] imm16  = instr_i[15:0];

// =====================================
// ����椸�]Decoder�^
// =====================================
Decoder DEC(
    .instr_op_i(opcode),
    .RegWrite_o(RegWrite_o),
    .MemtoReg_o(MemtoReg_o),
    .MemRead_o(MemRead_o),
    .MemWrite_o(MemWrite_o),
    .ALUSrc_o(ALUSrc_o),
    .ALUOp_o(ALUOp_o),
    .Branch_o(Branch_o)  
);

// =====================================
// Register File�]Ū�� rs�Brt�^
// =====================================
Reg_File RF(
    .clk      (clk),
    .rst      (rst),

    .RSaddr_i   (rs),
    .RTaddr_i   (rt),

    // ===== �g�^���q���g�J =====
    .RDaddr_i   (WB_WriteAddr_i),
    .RDdata_i   (WB_WriteData_i),
    .RegWrite_i (WB_RegWrite_i),

    // ===== ��X =====
    .RSdata_o   (rs_data_o),
    .RTdata_o   (rt_data_o)
);

// =====================================
// Sign Extend (branch address or immediate)
// =====================================
Sign_Extend SE(
    .data_i(imm16),
    .data_o(imm_o)
);

// =====================================
// Branch �P�_ (rs == rt ?)
// =====================================
assign Zero_o = (rs_data_o == rt_data_o);

// =====================================
// Branch Target Address
// PC + 4 + (imm << 2)
// =====================================
assign branch_target_o = pc_plus4_i + (imm_o << 2);

// =====================================
// ��X��}��T�� ID/EX
// =====================================
assign funct_o   = funct;
assign rs_addr_o = rs;
assign rt_addr_o = rt;
assign rd_addr_o = rd;

endmodule



