module ID_EX(
    input    clk,
    input    rst, 
    input ID_EX_Flush,      // hazard unit ����G1=�M��(ID/EX���JNOP), 0=���`��s
// Cycle 1: lw �b ID ���q
//          - Hazard Unit ������G�U�@���O�n�� lw �����G
//          - �o�X�H���GIF_ID_Write=0, PC_Write=0, ID_EX_Flush=0
         
// Cycle 2: lw �i EX�A�᭱���O�u�d�b IF/ID�v
//          - IF/ID ����s�]IF_ID_Write=0�^
//          - PC ���ʡ]PC_Write=0�^
//          - ID_EX �O����ȡ]ID_EX_Flush=0�A���`��s lw�^
//          - �᭱���O�٦b IF ���q�A�S�i ID
         
// Cycle 3: lw �i MEM�]���ɵ��G�i��X�ӤF�^
//          - �᭱���O�ש�i ID
//          - �Ϋe�X���� lw ���G�A�קK�A�d�@��

    // Control signals
    input RegWrite_i, MemtoReg_i, MemRead_i, MemWrite_i,
    // �O�_���\�⵲�G�g�^ Register File (R-type, lw, immmediate)
    // WB ���q�� mux ���� �Ӧ۰O�����٬O ALU (ALU(0) / Memory(1, lw))
    // �O����O�_�n���uŪ���v�ʧ@ (lw(1) / sw, R-type(0))
    // �O����O�_�n���u�g�J�v�ʧ@ (sw(1) / lw, R-type(0))
    input [1:0] ALUOp_i,                               // ALU control signals
    input ALUSrc_i,                                    // �M�w ALU ���ĤG�ӹB�⤸�Ӧۭ��� rt(0)/imm(1)

    // Data
    input [31:0] rs_i, rt_i, imm_i,                  // rs, rt, sign extended immediate
    input [5:0]  funct_i,                            // �P ALUOp �@�_�M�w ALU ����H��
    input [4:0]  rs_addr_i, rt_addr_i, rd_addr_i,    // �U���|���u

    // Outputs
    output reg RegWrite_o, MemtoReg_o, MemRead_o, MemWrite_o,
    output reg [1:0] ALUOp_o,
    output reg ALUSrc_o,

    output reg [31:0] rs_o, rt_o, imm_o,
    output reg [5:0]  funct_o,
    output reg [4:0]  rs_addr_o, rt_addr_o, rd_addr_o
);

always @(posedge clk or posedge rst) begin
    if (rst || ID_EX_Flush) begin
        {RegWrite_o, MemtoReg_o, MemRead_o, MemWrite_o} <= 0;
        ALUOp_o    <= 0;
        ALUSrc_o   <= 0;
        funct_o    <= 0;
        rs_o       <= 0;
        rt_o       <= 0;
        imm_o      <= 0;
        rs_addr_o  <= 0;
        rt_addr_o  <= 0;
        rd_addr_o  <= 0;
    end else begin
        RegWrite_o <= RegWrite_i;
        MemtoReg_o <= MemtoReg_i;
        MemRead_o  <= MemRead_i;
        MemWrite_o <= MemWrite_i;
        ALUOp_o    <= ALUOp_i;
        ALUSrc_o   <= ALUSrc_i;

        funct_o    <= funct_i;
        rs_o       <= rs_i;
        rt_o       <= rt_i;
        imm_o      <= imm_i;
        rs_addr_o  <= rs_addr_i;
        rt_addr_o  <= rt_addr_i;
        rd_addr_o  <= rd_addr_i;
    end
end

endmodule
