// =====================================
// WB Stage (Write Back)
// �t�d�G
//   - �ھ� MemtoReg �M�w�n�g�^ ALU ���G or Memory data
//   - �N���G��X�� Register File
// =====================================

module WB(
    // ===== MEM/WB pipeline inputs =====
    input         RegWrite_i,       // �O�_�n�g�^ RF
    input         MemtoReg_i,       // 1 = Memory data, 0 = ALU result
    input  [31:0] read_data_i,      // lw ���
    input  [31:0] ALU_result_i,     // R-type/addi/sw/lw �� ALU result
    input  [4:0]  dest_reg_i,       // �̲׭n�g�^�� register index

    // ===== outputs to Register File =====
    output        WB_RegWrite_o,    // �� RF ���g�J enable
    output [4:0]  WB_WriteAddr_o,   // �g�J���Ȧs���s��
    output [31:0] WB_WriteData_o    // �g�J�����
);

//
// =====================================
// 1. MemtoReg MUX
// =====================================
// �M�w�n�g�^���Ӹ��
assign WB_WriteData_o = (MemtoReg_i) ? read_data_i : ALU_result_i;      // to ALU mux and RF

//
// =====================================
// 2. �^�ǵ� Register File ������
// =====================================
assign WB_RegWrite_o  = RegWrite_i;    // �O�_�n�g�^, to forwarding unit and RF
assign WB_WriteAddr_o = dest_reg_i;    // �g�^���ӼȦs�� to forwarding unit and RF

endmodule
