module Instr_Memory(
    input  [31:0] addr_i,
    output [31:0] instr_o
);

reg [31:0] memory [0:255];  // 256 words (each 32-bit), �@ 1 KB ���O�O����

// ----------------------
// �q�ɮ׸��J���O
// ----------------------
initial begin
    // �N instruction.txt ���C�@�� HEX �̧Ǹ��J�� memory[0], memory[1], ...
    // �� 0 �� �� memory[0]
    // �� 1 �� �� memory[1]
    // �� N �� �� memory[N]
    $readmemb("instruction.txt", memory);
end

// ----------------------
// ���OŪ���]�ϥ� word addressing�^
// ----------------------
assign instr_o = memory[addr_i[31:2]];  
// �]�� MIPS ���O�O 4 bytes(32-bit)�APC �C���W�[ 4�C
// addr_i[31:2] ����� byte address �k�� 2�A�ন word index�C
// PC = 0 �� index=0
// PC = 4 �� index=1
// PC = 8 �� index=2

endmodule