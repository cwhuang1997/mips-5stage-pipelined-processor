// =====================================
// IF Stage (Instruction Fetch)
// �t�d�G
//   1. ���o PC
//   2. �q���O�O������X instr
//   3. �p�� PC + 4
//   4. ��X�� IF/ID pipeline register
// =====================================

module IF(
    input         clk,
    input         rst,
    input         PC_Write,        // hazard unit�G0 = stall ����s PC

    // ===== �Ӧ� ID stage �� branch �P�_ =====
    input         Branch_i,            // beq ���O�H
    input         Zero_i,              // rs == rt ?
    input  [31:0] branch_target_i,     // branch target address

    output [31:0] instr_o,         // �q IMEM ���X�����O
    output [31:0] pc_plus4_o,       // PC + 4 �� IF/ID


    output branch_taken_o
);


reg  [31:0] pc_reg;

// =====================================
// Branch �M���]PC ��ܾ��^
// branch_taken = Branch AND Zero
// =====================================
wire branch_taken = Branch_i & Zero_i;
assign branch_taken_o = branch_taken;

wire [31:0] pc_next = (branch_taken) ?
                      branch_target_i :   // branch �R�� �� ����ؼ�
                      pc_reg + 32'd4;     // otherwise �� PC + 4

// ===============================
// Program Counter (���ة󥻼Ҳ�)
// ===============================
always @(posedge clk or posedge rst) begin
    if (rst)
        pc_reg <= 32'b0;
    else if (PC_Write)
        pc_reg <= pc_next;   // ���`��s PC
    // else: PC_Write = 0 �� stall �� PC ����
end

// ===============================
// Instruction Memory
// ===============================
Instr_Memory IMEM(
    .addr_i(pc_reg),
    .instr_o(instr_o)
);

// ===============================
// PC + 4 �[�k��
// ===============================
assign pc_plus4_o = pc_reg + 32'd4;

endmodule
