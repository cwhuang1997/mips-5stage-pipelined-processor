// ===============================================
// Forwarding Unit
// �M�w EX ���q�ݭn�q���̨��B�⤸�G���` / EX/MEM / MEM/WB
// ===============================================
module Forwarding_Unit(

    // ===== �Ӧ� ID/EX (�{����O�ϥΪ��Ȧs��) =====
    input  [4:0] ID_EX_rs,          // EX ���q�i�Ӫ�rs �h��Ӧ��S����᭱�n�g�^���@��
    input  [4:0] ID_EX_rt,          // EX ���q�i�Ӫ�rt �h��Ӧ��S����᭱�n�g�^���@��

    // ===== �Ӧ� EX/MEM (�W�@�����O) =====
    input        EX_MEM_RegWrite,
    input  [4:0] EX_MEM_rd,          // EX/MEM dest register

    // ===== �Ӧ� MEM/WB (�A�W�@�����O) =====
    input        MEM_WB_RegWrite,
    input  [4:0] MEM_WB_rd,          // MEM/WB dest register

    // ===== Forwarding outputs =====
    output reg [1:0] ForwardA,
    output reg [1:0] ForwardB
);

always @(*) begin
    // �w�]�� forward
    ForwardA = 2'b00;
    ForwardB = 2'b00;

    // ====================================
    // Forward A (src1)
    // ====================================
    // EX hazard�GEX/MEM �� EX
    if (EX_MEM_RegWrite &&
        (EX_MEM_rd != 0) &&
        (EX_MEM_rd == ID_EX_rs)) begin
        ForwardA = 2'b10;
    end
    // MEM hazard�GMEM/WB �� EX
    else if (MEM_WB_RegWrite &&
             (MEM_WB_rd != 0) &&
             (MEM_WB_rd == ID_EX_rs)) begin
        ForwardA = 2'b01;
    end

    // ====================================
    // Forward B (src2)
    // ====================================
    if (EX_MEM_RegWrite &&
        (EX_MEM_rd != 0) &&
        (EX_MEM_rd == ID_EX_rt)) begin
        ForwardB = 2'b10;
    end
    else if (MEM_WB_RegWrite &&
             (MEM_WB_rd != 0) &&
             (MEM_WB_rd == ID_EX_rt)) begin
        ForwardB = 2'b01;
    end
end

endmodule
